module main

pub interface Form {
	color Volor
	hit(Vay) ?Vector3
}
