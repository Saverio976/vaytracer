module vtc

import gg

pub struct Material {
	color     gg.Color
	ambient   f64
	diffuse   f64
	specular  f64
	shininess f64
}
