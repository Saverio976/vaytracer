module vtc

pub struct Color {
pub mut:
	r u8
	g u8
	b u8
	a u8 = 255
}
