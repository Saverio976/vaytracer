module vtc

import math.vec

pub struct Vay {
pub mut:
	origin    vec.Vec3[f64]
	direction vec.Vec3[f64]
}
