module main

pub struct Volor {
pub:
	r u8
	g u8
	b u8
	a u8
}
