module vtc

pub struct Material {
	color     Color
	ambient   f64
	diffuse   f64
	specular  f64
	shininess f64
}
